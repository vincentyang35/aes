`ifndef AES_PKG_SV
`define AES_PKG_SV
package aes_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "aes_tx.sv"
  `include "aes_config.sv"
  `include "aes_driver.sv"
  `include "aes_monitor.sv"
  `include "aes_sequencer.sv"
  `include "aes_coverage.sv"
  `include "aes_agent.sv"
  `include "sequences/aes_seq_lib.sv"
  `include "sequences/aes_top_seq_lib.sv"
endpackage : aes_pkg

`endif  // AES_PKG_SV
