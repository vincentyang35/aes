`ifndef AES_SEQUENCER_SV
`define AES_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(aes_tx) aes_sequencer_t;


`endif // AES_SEQUENCER_SV
